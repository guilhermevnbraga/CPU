module cpu 
	(output reg [7:0] address,
	 output reg [7:0] to_memory
	 output reg write,
	 input wire [7:0] from_memory, 
     input wire clk, reset);
             
  	// Complement the module

endmodule